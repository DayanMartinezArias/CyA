module puerta_and3 (output wire y, input wire a,b,c);
  assign y = a & b & c;
endmodule